`timescale 1ns / 1ps
/*
`define DATA_X 28
`define DATA_Y 28
`define DATA_SIZE 32
`define WEIGHT_X 5
`define WEIGHT_Y 5
`define WEIGHT_SIZE 32
`define WEIGHT_WIDTH 32
`define CONV_X 24
`define CONV_Y 24
`define CONV_SIZE 69
`define RELU_X 24
`define RELU_Y 24
`define RELU_DATA_WIDTH 69
`define POOL_X 12
`define POOL_Y 12
`define STRIDE 2
*/
module simpleCNN (
	input wire clk,    // Clock
	input wire rst,  	// Asynchronous reset active high
	input wire enable,
	output reg [3:0] result,
	output reg [15:0] count,
	output wire signed [112:0] prob_0,
	output wire signed [112:0] prob_1,
	output wire signed [112:0] prob_2,
	output wire signed [112:0] prob_3,
	output wire signed [112:0] prob_4,
	output wire signed [112:0] prob_5,
	output wire signed [112:0] prob_6,
	output wire signed [112:0] prob_7,
	output wire signed [112:0] prob_8,
	output wire signed [112:0] prob_9,
	output wire fc_done
);
	reg signed [112:0] prob [9:0];
	integer i,j;
// conv_layer
	wire signed [68:0] conv_result_1;
	wire signed [68:0] conv_result_2;
	wire signed [68:0] conv_result_3;
	wire signed [68:0] conv_result_4;
	wire signed [68:0] conv_result_5;
	wire signed [68:0] conv_result_6;
	wire signed [68:0] conv_result_7;
	wire signed [68:0] conv_result_8;
// relu_layer
	wire signed [68:0] relu_result_1;
	wire signed [68:0] relu_result_2;
	wire signed [68:0] relu_result_3;
	wire signed [68:0] relu_result_4;
	wire signed [68:0] relu_result_5;
	wire signed [68:0] relu_result_6;
	wire signed [68:0] relu_result_7;
	wire signed [68:0] relu_result_8;
// pool_layer
	wire signed [68:0] pool_result_1;
	wire signed [68:0] pool_result_2;
	wire signed [68:0] pool_result_3;
	wire signed [68:0] pool_result_4;
	wire signed [68:0] pool_result_5;
	wire signed [68:0] pool_result_6;
	wire signed [68:0] pool_result_7;
	wire signed [68:0] pool_result_8;
// fc_layer
/*
	wire signed [112:0] prob_0;
	wire signed [112:0] prob_1;
	wire signed [112:0] prob_2;
	wire signed [112:0] prob_3;
	wire signed [112:0] prob_4;
	wire signed [112:0] prob_5;
	wire signed [112:0] prob_6;
	wire signed [112:0] prob_7;
	wire signed [112:0] prob_8;
	wire signed [112:0] prob_9;
	wire fc_done;
*/
	reg [4:0] count_x, relu_count_x;
	reg [4:0] count_y, relu_count_y;
	//reg [15:0] count;
	wire signed [31:0] data [0:27][0:27];
	reg data_read_done;
	reg signed [68:0] relu [7:0][575:0];
	reg signed [68:0] relu_1 [23:0][23:0];
	reg signed [68:0] relu_2 [23:0][23:0];
	reg signed [68:0] relu_3 [23:0][23:0];
	reg signed [68:0] relu_4 [23:0][23:0];
	reg signed [68:0] relu_5 [23:0][23:0];
	reg signed [68:0] relu_6 [23:0][23:0];
	reg signed [68:0] relu_7 [23:0][23:0];
	reg signed [68:0] relu_8 [23:0][23:0];
	reg signed [68:0] pool [7:0][143:0];
	reg signed [31:0] data_00;
	reg signed [31:0] data_01;
	reg signed [31:0] data_02;
	reg signed [31:0] data_03;
	reg signed [31:0] data_04;
	reg signed [31:0] data_10;
	reg signed [31:0] data_11;
	reg signed [31:0] data_12;
	reg signed [31:0] data_13;
	reg signed [31:0] data_14;
	reg signed [31:0] data_20;
	reg signed [31:0] data_21;
	reg signed [31:0] data_22;
	reg signed [31:0] data_23;
	reg signed [31:0] data_24;
	reg signed [31:0] data_30;
	reg signed [31:0] data_31;
	reg signed [31:0] data_32;
	reg signed [31:0] data_33;
	reg signed [31:0] data_34;
	reg signed [31:0] data_40;
	reg signed [31:0] data_41;
	reg signed [31:0] data_42;
	reg signed [31:0] data_43;
	reg signed [31:0] data_44;
	reg signed [68:0] pool_0_00;
	reg signed [68:0] pool_0_01;
	reg signed [68:0] pool_0_10;
	reg signed [68:0] pool_0_11;
	reg signed [68:0] pool_1_00;
	reg signed [68:0] pool_1_01;
	reg signed [68:0] pool_1_10;
	reg signed [68:0] pool_1_11;
	reg signed [68:0] pool_2_00;
	reg signed [68:0] pool_2_01;
	reg signed [68:0] pool_2_10;
	reg signed [68:0] pool_2_11;
	reg signed [68:0] pool_3_00;
	reg signed [68:0] pool_3_01;
	reg signed [68:0] pool_3_10;
	reg signed [68:0] pool_3_11;
	reg signed [68:0] pool_4_00;
	reg signed [68:0] pool_4_01;
	reg signed [68:0] pool_4_10;
	reg signed [68:0] pool_4_11;
	reg signed [68:0] pool_5_00;
	reg signed [68:0] pool_5_01;
	reg signed [68:0] pool_5_10;
	reg signed [68:0] pool_5_11;
	reg signed [68:0] pool_6_00;
	reg signed [68:0] pool_6_01;
	reg signed [68:0] pool_6_10;
	reg signed [68:0] pool_6_11;
	reg signed [68:0] pool_7_00;
	reg signed [68:0] pool_7_01;
	reg signed [68:0] pool_7_10;
	reg signed [68:0] pool_7_11;

assign data[0][0] = 32'b00000000001101000011010000110100;
assign data[0][1] = 32'b00000000000000110101100010101110;
assign data[0][2] = 32'b00000000000000000000000000000000;
assign data[0][3] = 32'b00000000000000000000000000000000;
assign data[0][4] = 32'b00000000000000000000000000000000;
assign data[0][5] = 32'b00000000000000000000000000000000;
assign data[0][6] = 32'b00000000000000000000000000000000;
assign data[0][7] = 32'b00000000000000000000000000000000;
assign data[0][8] = 32'b00000000000000000000000000000000;
assign data[0][9] = 32'b00000000000000000000000000000000;
assign data[0][10] = 32'b00000000000000000000000000000000;
assign data[0][11] = 32'b00000000000000000000000000000000;
assign data[0][12] = 32'b00000000000000000000000000000000;
assign data[0][13] = 32'b00000000000000000000000000000000;
assign data[0][14] = 32'b00000000000000000000000000000000;
assign data[0][15] = 32'b00000000000000000000000000000000;
assign data[0][16] = 32'b00000000000000000000000000000000;
assign data[0][17] = 32'b00000000000000000000000000000000;
assign data[0][18] = 32'b00000000000000000000000000000000;
assign data[0][19] = 32'b00000000000000000000000000000000;
assign data[0][20] = 32'b00000000000000000000000000000000;
assign data[0][21] = 32'b00000000000000000000000000000000;
assign data[0][22] = 32'b00000000000000000000000000000000;
assign data[0][23] = 32'b00000000000000000000000000000000;
assign data[0][24] = 32'b00000000000000000000000000000000;
assign data[0][25] = 32'b00000000000000000000000000000000;
assign data[0][26] = 32'b00000000000000000000000000000000;
assign data[0][27] = 32'b00000000000000000000000000000000;
assign data[1][0] = 32'b00000000000000000000000000000000;
assign data[1][1] = 32'b00000000000000000000000000000000;
assign data[1][2] = 32'b00000000000000000000000000000000;
assign data[1][3] = 32'b00000000000000000000000000000000;
assign data[1][4] = 32'b00000000000000000000000000000000;
assign data[1][5] = 32'b00000000000000000000000000000000;
assign data[1][6] = 32'b00000000000000000000000000000000;
assign data[1][7] = 32'b00000000000000000000000000000000;
assign data[1][8] = 32'b00000000000000000000000000000000;
assign data[1][9] = 32'b00000000000000000000000000000000;
assign data[1][10] = 32'b00000000000000000000000000000000;
assign data[1][11] = 32'b00000000000000000000000000000000;
assign data[1][12] = 32'b00000000000000000000000000000000;
assign data[1][13] = 32'b00000000000000000000000000000000;
assign data[1][14] = 32'b00000000000000000000000000000000;
assign data[1][15] = 32'b00000000000000000000000000000000;
assign data[1][16] = 32'b00000000000000000000000000000000;
assign data[1][17] = 32'b00000000000000000000000000000000;
assign data[1][18] = 32'b00000000000000000000000000000000;
assign data[1][19] = 32'b00000000000000000000000000000000;
assign data[1][20] = 32'b00000000000000000000000000000000;
assign data[1][21] = 32'b00000000000000000000000000000000;
assign data[1][22] = 32'b00000000000000000000000000000000;
assign data[1][23] = 32'b00000000000000000000000000000000;
assign data[1][24] = 32'b00000000000000000000000000000000;
assign data[1][25] = 32'b00000000000000000000000000000000;
assign data[1][26] = 32'b00000000000000000000000000000000;
assign data[1][27] = 32'b00000000000000000000000000000000;
assign data[2][0] = 32'b00000000000000000000000000000000;
assign data[2][1] = 32'b00000000000000000000000000000000;
assign data[2][2] = 32'b00000000000000000000000000000000;
assign data[2][3] = 32'b00000000000000000000000000000000;
assign data[2][4] = 32'b00000000000000000000000000000000;
assign data[2][5] = 32'b00000000000000000000000000000000;
assign data[2][6] = 32'b00000000000000000000000000000000;
assign data[2][7] = 32'b00000000000000000000000000000000;
assign data[2][8] = 32'b00000000000000000000000000000000;
assign data[2][9] = 32'b00000000000000000000000000000000;
assign data[2][10] = 32'b00000000000000000000000000000000;
assign data[2][11] = 32'b00000000000000000000000000000000;
assign data[2][12] = 32'b00000000000000000000000000000000;
assign data[2][13] = 32'b00000000000000000000000000000000;
assign data[2][14] = 32'b00000000000000000000000000000000;
assign data[2][15] = 32'b00000000000000000000000000000000;
assign data[2][16] = 32'b00000000000000000000000000000000;
assign data[2][17] = 32'b00000000000000000000000000000000;
assign data[2][18] = 32'b00000000000000000000000000000000;
assign data[2][19] = 32'b00000000000000000000000000000000;
assign data[2][20] = 32'b00000000000000000000000000000000;
assign data[2][21] = 32'b00000000000000000000000000000000;
assign data[2][22] = 32'b00000000000000000000000000000000;
assign data[2][23] = 32'b00000000000000000000000000000000;
assign data[2][24] = 32'b00000000000000000000000000000000;
assign data[2][25] = 32'b00000000000000000000000000000000;
assign data[2][26] = 32'b00000000000000000000000000000000;
assign data[2][27] = 32'b00000000000000000000000000000000;
assign data[3][0] = 32'b00000000000000000000000000000000;
assign data[3][1] = 32'b00000000000000000000000000000000;
assign data[3][2] = 32'b00000000000000000000000000000000;
assign data[3][3] = 32'b00000000000000000000000000000000;
assign data[3][4] = 32'b00000000000000000000000000000000;
assign data[3][5] = 32'b00000000000000000000000000000000;
assign data[3][6] = 32'b00000000000000000000000000000000;
assign data[3][7] = 32'b00000000000000000000000000000000;
assign data[3][8] = 32'b00000000000000000000000000000000;
assign data[3][9] = 32'b00000000000000000000000000000000;
assign data[3][10] = 32'b00000000000000000000000000000000;
assign data[3][11] = 32'b00000000000000000000000000000000;
assign data[3][12] = 32'b00000000000000000000000000000000;
assign data[3][13] = 32'b00000000000000000000000000000000;
assign data[3][14] = 32'b00000000000000000000000000000000;
assign data[3][15] = 32'b00000000000000000000000000000000;
assign data[3][16] = 32'b00000000000000000000000000000000;
assign data[3][17] = 32'b00000000000000000000000000000000;
assign data[3][18] = 32'b00000000000000000000000000000000;
assign data[3][19] = 32'b00000000000000000000000000000000;
assign data[3][20] = 32'b00000000000000000000000000000000;
assign data[3][21] = 32'b00000000000000000000000000000000;
assign data[3][22] = 32'b00000000000000000000000000000000;
assign data[3][23] = 32'b00000000000000000000000000000000;
assign data[3][24] = 32'b00000000000000000000000000000000;
assign data[3][25] = 32'b00000000000000000000000000000000;
assign data[3][26] = 32'b00000000000000000000000000000000;
assign data[3][27] = 32'b00000000000000000000000000000000;
assign data[4][0] = 32'b00000000000000000000000000000000;
assign data[4][1] = 32'b00000000000000000000000000000000;
assign data[4][2] = 32'b00000000000000000000000000000000;
assign data[4][3] = 32'b00000000000000000000000000000000;
assign data[4][4] = 32'b00000000000000000000000000000000;
assign data[4][5] = 32'b00000000000000000000000000000000;
assign data[4][6] = 32'b00000000000000000000000000000000;
assign data[4][7] = 32'b00000000000000000000000000000000;
assign data[4][8] = 32'b00000000000000000000000000000000;
assign data[4][9] = 32'b00000000000000000000000000000000;
assign data[4][10] = 32'b00000000000000000000000000000000;
assign data[4][11] = 32'b00000000000000000000000000000000;
assign data[4][12] = 32'b00000000000000000000000000000000;
assign data[4][13] = 32'b00000000000000000000000000000000;
assign data[4][14] = 32'b00000000000000000000000000000000;
assign data[4][15] = 32'b00000000000000000000000000000000;
assign data[4][16] = 32'b00000000000000000000000000000000;
assign data[4][17] = 32'b00000000000000000000000000000000;
assign data[4][18] = 32'b00000000000000000000000000000000;
assign data[4][19] = 32'b00000000000000000000000000000000;
assign data[4][20] = 32'b00000000000000000000000000000000;
assign data[4][21] = 32'b00000000000000000000000000000000;
assign data[4][22] = 32'b00000000000000000000000000000000;
assign data[4][23] = 32'b00000000000000000000000000000000;
assign data[4][24] = 32'b00000000000000000000000000000000;
assign data[4][25] = 32'b00000000000000000000000000000000;
assign data[4][26] = 32'b00000000000000000000000000000000;
assign data[4][27] = 32'b00000000000000000000000000000000;
assign data[5][0] = 32'b00000000000000000000000000000000;
assign data[5][1] = 32'b00000000000000000000000000000000;
assign data[5][2] = 32'b00000000000000000000000000000000;
assign data[5][3] = 32'b00000000000000000000000000000000;
assign data[5][4] = 32'b00000000000000000000000000000000;
assign data[5][5] = 32'b00000000000000000000000000000000;
assign data[5][6] = 32'b00000000000000000000000000000000;
assign data[5][7] = 32'b00000000000000000000000000000000;
assign data[5][8] = 32'b00000000000000000000000000000000;
assign data[5][9] = 32'b00000000000000000000000000000000;
assign data[5][10] = 32'b00000000000000000000000000000000;
assign data[5][11] = 32'b00000000000000000000000000000000;
assign data[5][12] = 32'b00000000000000000000000000000000;
assign data[5][13] = 32'b00000000000000000000000000000000;
assign data[5][14] = 32'b00000000000000000000000000000000;
assign data[5][15] = 32'b00000000000000000000000000000000;
assign data[5][16] = 32'b00000000000000000000000000000000;
assign data[5][17] = 32'b00000000000000000000000000000000;
assign data[5][18] = 32'b00000000000000000000000000000000;
assign data[5][19] = 32'b00000000000000000000000000000000;
assign data[5][20] = 32'b00000000000000000000000000000000;
assign data[5][21] = 32'b00000000000000000000000000000000;
assign data[5][22] = 32'b00000000000000000000000000000000;
assign data[5][23] = 32'b00000000000000000000000000000000;
assign data[5][24] = 32'b00000000000000000000000000000000;
assign data[5][25] = 32'b00000000000000000000000000000000;
assign data[5][26] = 32'b00000000000000000000000000000000;
assign data[5][27] = 32'b00000000000000000000000000000000;
assign data[6][0] = 32'b00000000000000000000000000000000;
assign data[6][1] = 32'b00000000000000000000000000000000;
assign data[6][2] = 32'b00000000000000000000000000000000;
assign data[6][3] = 32'b00000000000000000000000000000000;
assign data[6][4] = 32'b00000000000000000000000000000000;
assign data[6][5] = 32'b00000000000000000000000000000000;
assign data[6][6] = 32'b00000000000000000000000000000000;
assign data[6][7] = 32'b00000000000000010101011010101100;
assign data[6][8] = 32'b00000000000010100000101000001010;
assign data[6][9] = 32'b00000000000011100000111000001110;
assign data[6][10] = 32'b00000000000001100000011000000110;
assign data[6][11] = 32'b00000000000000001010101101010110;
assign data[6][12] = 32'b00000000000000000000000000000000;
assign data[6][13] = 32'b00000000000000000000000000000000;
assign data[6][14] = 32'b00000000000000000000000000000000;
assign data[6][15] = 32'b00000000000000000000000000000000;
assign data[6][16] = 32'b00000000000000000000000000000000;
assign data[6][17] = 32'b00000000000000000000000000000000;
assign data[6][18] = 32'b00000000000000000000000000000000;
assign data[6][19] = 32'b00000000000000000000000000000000;
assign data[6][20] = 32'b00000000000000000000000000000000;
assign data[6][21] = 32'b00000000000000000000000000000000;
assign data[6][22] = 32'b00000000000000000000000000000000;
assign data[6][23] = 32'b00000000000000000000000000000000;
assign data[6][24] = 32'b00000000000000000000000000000000;
assign data[6][25] = 32'b00000000000000000000000000000000;
assign data[6][26] = 32'b00000000000000000000000000000000;
assign data[6][27] = 32'b00000000000000000000000000000000;
assign data[7][0] = 32'b00000000000000000000000000000000;
assign data[7][1] = 32'b00000000000000000000000000000000;
assign data[7][2] = 32'b00000000000000000000000000000000;
assign data[7][3] = 32'b00000000000000000000000000000000;
assign data[7][4] = 32'b00000000000000000000000000000000;
assign data[7][5] = 32'b00000000000000000000000000000000;
assign data[7][6] = 32'b00000000000000000000000000000000;
assign data[7][7] = 32'b00000000000011101011100101100100;
assign data[7][8] = 32'b00000000010101011010101100000001;
assign data[7][9] = 32'b00000000011110100010010011010000;
assign data[7][10] = 32'b00000000011011111100010100011011;
assign data[7][11] = 32'b00000000010111000000011010110010;
assign data[7][12] = 32'b00000000010011001010000111111000;
assign data[7][13] = 32'b00000000001111101110100110010100;
assign data[7][14] = 32'b00000000001100101101110110001000;
assign data[7][15] = 32'b00000000001001000111100111001111;
assign data[7][16] = 32'b00000000000111011100100001110011;
assign data[7][17] = 32'b00000000000100100110011110111101;
assign data[7][18] = 32'b00000000000001010000010100000101;
assign data[7][19] = 32'b00000000000000000101010110101011;
assign data[7][20] = 32'b00000000000000000000000000000000;
assign data[7][21] = 32'b00000000000000000000000000000000;
assign data[7][22] = 32'b00000000000000000000000000000000;
assign data[7][23] = 32'b00000000000000000000000000000000;
assign data[7][24] = 32'b00000000000000000000000000000000;
assign data[7][25] = 32'b00000000000000000000000000000000;
assign data[7][26] = 32'b00000000000000000000000000000000;
assign data[7][27] = 32'b00000000000000000000000000000000;
assign data[8][0] = 32'b00000000000000000000000000000000;
assign data[8][1] = 32'b00000000000000000000000000000000;
assign data[8][2] = 32'b00000000000000000000000000000000;
assign data[8][3] = 32'b00000000000000000000000000000000;
assign data[8][4] = 32'b00000000000000000000000000000000;
assign data[8][5] = 32'b00000000000000000000000000000000;
assign data[8][6] = 32'b00000000000000000000000000000000;
assign data[8][7] = 32'b00000000001100011000011011011100;
assign data[8][8] = 32'b00000000101001110101000111111101;
assign data[8][9] = 32'b00000000110111110011010010001010;
assign data[8][10] = 32'b00000000111001110011110010010010;
assign data[8][11] = 32'b00000000111000111000111000111001;
assign data[8][12] = 32'b00000000110101101101011011010111;
assign data[8][13] = 32'b00000000110001110001110001110010;
assign data[8][14] = 32'b00000000101101111011011110111000;
assign data[8][15] = 32'b00000000101001001010010010100101;
assign data[8][16] = 32'b00000000100110000100001011101110;
assign data[8][17] = 32'b00000000100001100011000011011100;
assign data[8][18] = 32'b00000000011001000110010001100101;
assign data[8][19] = 32'b00000000010010011111010010100000;
assign data[8][20] = 32'b00000000001110110011101100111011;
assign data[8][21] = 32'b00000000001000111100111001111001;
assign data[8][22] = 32'b00000000000010101011010101100000;
assign data[8][23] = 32'b00000000000000010000000100000001;
assign data[8][24] = 32'b00000000000000000000000000000000;
assign data[8][25] = 32'b00000000000000000000000000000000;
assign data[8][26] = 32'b00000000000000000000000000000000;
assign data[8][27] = 32'b00000000000000000000000000000000;
assign data[9][0] = 32'b00000000000000000000000000000000;
assign data[9][1] = 32'b00000000000000000000000000000000;
assign data[9][2] = 32'b00000000000000000000000000000000;
assign data[9][3] = 32'b00000000000000000000000000000000;
assign data[9][4] = 32'b00000000000000000000000000000000;
assign data[9][5] = 32'b00000000000000000000000000000000;
assign data[9][6] = 32'b00000000000000000000000000000000;
assign data[9][7] = 32'b00000000000001101011000101011100;
assign data[9][8] = 32'b00000000001110001110001110001110;
assign data[9][9] = 32'b00000000010101111010110100000011;
assign data[9][10] = 32'b00000000011001100001000010111100;
assign data[9][11] = 32'b00000000011111000010011011010010;
assign data[9][12] = 32'b00000000100100111110100100111111;
assign data[9][13] = 32'b00000000101010001111111001010100;
assign data[9][14] = 32'b00000000101110110001000001100110;
assign data[9][15] = 32'b00000000110010010111010000011111;
assign data[9][16] = 32'b00000000110101011101010111010110;
assign data[9][17] = 32'b00000000110111011101110111011110;
assign data[9][18] = 32'b00000000110110010010111010000100;
assign data[9][19] = 32'b00000000110011010010001001111000;
assign data[9][20] = 32'b00000000110000010110110000010111;
assign data[9][21] = 32'b00000000100100011001000110010010;
assign data[9][22] = 32'b00000000001110001000110111100011;
assign data[9][23] = 32'b00000000000001111011001001011101;
assign data[9][24] = 32'b00000000000000000000000000000000;
assign data[9][25] = 32'b00000000000000000000000000000000;
assign data[9][26] = 32'b00000000000000000000000000000000;
assign data[9][27] = 32'b00000000000000000000000000000000;
assign data[10][0] = 32'b00000000000000000000000000000000;
assign data[10][1] = 32'b00000000000000000000000000000000;
assign data[10][2] = 32'b00000000000000000000000000000000;
assign data[10][3] = 32'b00000000000000000000000000000000;
assign data[10][4] = 32'b00000000000000000000000000000000;
assign data[10][5] = 32'b00000000000000000000000000000000;
assign data[10][6] = 32'b00000000000000000000000000000000;
assign data[10][7] = 32'b00000000000000000000000000000000;
assign data[10][8] = 32'b00000000000000000000000000000000;
assign data[10][9] = 32'b00000000000000000000000000000000;
assign data[10][10] = 32'b00000000000000010101011010101100;
assign data[10][11] = 32'b00000000000011000000110000001100;
assign data[10][12] = 32'b00000000000110111100011001110001;
assign data[10][13] = 32'b00000000001010011101010001111111;
assign data[10][14] = 32'b00000000001101101110000110001100;
assign data[10][15] = 32'b00000000010000110100001101000100;
assign data[10][16] = 32'b00000000010100010101000101010010;
assign data[10][17] = 32'b00000000011010100110101001101011;
assign data[10][18] = 32'b00000000100001110011000111011101;
assign data[10][19] = 32'b00000000101100001011000010110001;
assign data[10][20] = 32'b00000000110100010111110000100111;
assign data[10][21] = 32'b00000000101100100101110100001000;
assign data[10][22] = 32'b00000000010011011010001011111001;
assign data[10][23] = 32'b00000000000011000110000110110111;
assign data[10][24] = 32'b00000000000000000000000000000000;
assign data[10][25] = 32'b00000000000000000000000000000000;
assign data[10][26] = 32'b00000000000000000000000000000000;
assign data[10][27] = 32'b00000000000000000000000000000000;
assign data[11][0] = 32'b00000000000000000000000000000000;
assign data[11][1] = 32'b00000000000000000000000000000000;
assign data[11][2] = 32'b00000000000000000000000000000000;
assign data[11][3] = 32'b00000000000000000000000000000000;
assign data[11][4] = 32'b00000000000000000000000000000000;
assign data[11][5] = 32'b00000000000000000000000000000000;
assign data[11][6] = 32'b00000000000000000000000000000000;
assign data[11][7] = 32'b00000000000000000000000000000000;
assign data[11][8] = 32'b00000000000000000000000000000000;
assign data[11][9] = 32'b00000000000000000000000000000000;
assign data[11][10] = 32'b00000000000000000000000000000000;
assign data[11][11] = 32'b00000000000000000000000000000000;
assign data[11][12] = 32'b00000000000000000000000000000000;
assign data[11][13] = 32'b00000000000000000000000000000000;
assign data[11][14] = 32'b00000000000000000000000000000000;
assign data[11][15] = 32'b00000000000000000000000000000000;
assign data[11][16] = 32'b00000000000000001010101101010110;
assign data[11][17] = 32'b00000000000001111011001001011101;
assign data[11][18] = 32'b00000000001110111110011010010001;
assign data[11][19] = 32'b00000000101001011111101101010001;
assign data[11][20] = 32'b00000000110101111000001000101101;
assign data[11][21] = 32'b00000000100111101111010001001010;
assign data[11][22] = 32'b00000000001101100011011000110110;
assign data[11][23] = 32'b00000000000001011011000001011011;
assign data[11][24] = 32'b00000000000000000000000000000000;
assign data[11][25] = 32'b00000000000000000000000000000000;
assign data[11][26] = 32'b00000000000000000000000000000000;
assign data[11][27] = 32'b00000000000000000000000000000000;
assign data[12][0] = 32'b00000000000000000000000000000000;
assign data[12][1] = 32'b00000000000000000000000000000000;
assign data[12][2] = 32'b00000000000000000000000000000000;
assign data[12][3] = 32'b00000000000000000000000000000000;
assign data[12][4] = 32'b00000000000000000000000000000000;
assign data[12][5] = 32'b00000000000000000000000000000000;
assign data[12][6] = 32'b00000000000000000000000000000000;
assign data[12][7] = 32'b00000000000000000000000000000000;
assign data[12][8] = 32'b00000000000000000000000000000000;
assign data[12][9] = 32'b00000000000000000000000000000000;
assign data[12][10] = 32'b00000000000000000000000000000000;
assign data[12][11] = 32'b00000000000000000000000000000000;
assign data[12][12] = 32'b00000000000000000000000000000000;
assign data[12][13] = 32'b00000000000000000000000000000000;
assign data[12][14] = 32'b00000000000000000000000000000000;
assign data[12][15] = 32'b00000000000000000000000000000000;
assign data[12][16] = 32'b00000000000000000000000000000000;
assign data[12][17] = 32'b00000000000011110110010010111010;
assign data[12][18] = 32'b00000000011011010110110101101110;
assign data[12][19] = 32'b00000000110001000001100101101111;
assign data[12][20] = 32'b00000000101011000101011100000010;
assign data[12][21] = 32'b00000000010001011111000010011100;
assign data[12][22] = 32'b00000000000010110110000010110110;
assign data[12][23] = 32'b00000000000000001010101101010110;
assign data[12][24] = 32'b00000000000000000000000000000000;
assign data[12][25] = 32'b00000000000000000000000000000000;
assign data[12][26] = 32'b00000000000000000000000000000000;
assign data[12][27] = 32'b00000000000000000000000000000000;
assign data[13][0] = 32'b00000000000000000000000000000000;
assign data[13][1] = 32'b00000000000000000000000000000000;
assign data[13][2] = 32'b00000000000000000000000000000000;
assign data[13][3] = 32'b00000000000000000000000000000000;
assign data[13][4] = 32'b00000000000000000000000000000000;
assign data[13][5] = 32'b00000000000000000000000000000000;
assign data[13][6] = 32'b00000000000000000000000000000000;
assign data[13][7] = 32'b00000000000000000000000000000000;
assign data[13][8] = 32'b00000000000000000000000000000000;
assign data[13][9] = 32'b00000000000000000000000000000000;
assign data[13][10] = 32'b00000000000000000000000000000000;
assign data[13][11] = 32'b00000000000000000000000000000000;
assign data[13][12] = 32'b00000000000000000000000000000000;
assign data[13][13] = 32'b00000000000000000000000000000000;
assign data[13][14] = 32'b00000000000000000000000000000000;
assign data[13][15] = 32'b00000000000000000000000000000000;
assign data[13][16] = 32'b00000000000000001010101101010110;
assign data[13][17] = 32'b00000000001101011110000010001011;
assign data[13][18] = 32'b00000000101001010100111111111011;
assign data[13][19] = 32'b00000000101111100110100100010100;
assign data[13][20] = 32'b00000000011000000000101010110110;
assign data[13][21] = 32'b00000000000100100110011110111101;
assign data[13][22] = 32'b00000000000000000101010110101011;
assign data[13][23] = 32'b00000000000000000000000000000000;
assign data[13][24] = 32'b00000000000000000000000000000000;
assign data[13][25] = 32'b00000000000000000000000000000000;
assign data[13][26] = 32'b00000000000000000000000000000000;
assign data[13][27] = 32'b00000000000000000000000000000000;
assign data[14][0] = 32'b00000000000000000000000000000000;
assign data[14][1] = 32'b00000000000000000000000000000000;
assign data[14][2] = 32'b00000000000000000000000000000000;
assign data[14][3] = 32'b00000000000000000000000000000000;
assign data[14][4] = 32'b00000000000000000000000000000000;
assign data[14][5] = 32'b00000000000000000000000000000000;
assign data[14][6] = 32'b00000000000000000000000000000000;
assign data[14][7] = 32'b00000000000000000000000000000000;
assign data[14][8] = 32'b00000000000000000000000000000000;
assign data[14][9] = 32'b00000000000000000000000000000000;
assign data[14][10] = 32'b00000000000000000000000000000000;
assign data[14][11] = 32'b00000000000000000000000000000000;
assign data[14][12] = 32'b00000000000000000000000000000000;
assign data[14][13] = 32'b00000000000000000000000000000000;
assign data[14][14] = 32'b00000000000000000000000000000000;
assign data[14][15] = 32'b00000000000000000000000000000000;
assign data[14][16] = 32'b00000000000010110110000010110110;
assign data[14][17] = 32'b00000000011000100000110010111000;
assign data[14][18] = 32'b00000000101111101011111010111111;
assign data[14][19] = 32'b00000000100101010011111111101011;
assign data[14][20] = 32'b00000000001011001000000111010111;
assign data[14][21] = 32'b00000000000000110000001100000011;
assign data[14][22] = 32'b00000000000000000000000000000000;
assign data[14][23] = 32'b00000000000000000000000000000000;
assign data[14][24] = 32'b00000000000000000000000000000000;
assign data[14][25] = 32'b00000000000000000000000000000000;
assign data[14][26] = 32'b00000000000000000000000000000000;
assign data[14][27] = 32'b00000000000000000000000000000000;
assign data[15][0] = 32'b00000000000000000000000000000000;
assign data[15][1] = 32'b00000000000000000000000000000000;
assign data[15][2] = 32'b00000000000000000000000000000000;
assign data[15][3] = 32'b00000000000000000000000000000000;
assign data[15][4] = 32'b00000000000000000000000000000000;
assign data[15][5] = 32'b00000000000000000000000000000000;
assign data[15][6] = 32'b00000000000000000000000000000000;
assign data[15][7] = 32'b00000000000000000000000000000000;
assign data[15][8] = 32'b00000000000000000000000000000000;
assign data[15][9] = 32'b00000000000000000000000000000000;
assign data[15][10] = 32'b00000000000000000000000000000000;
assign data[15][11] = 32'b00000000000000000000000000000000;
assign data[15][12] = 32'b00000000000000000000000000000000;
assign data[15][13] = 32'b00000000000000000000000000000000;
assign data[15][14] = 32'b00000000000000000000000000000000;
assign data[15][15] = 32'b00000000000000010101011010101100;
assign data[15][16] = 32'b00000000001101001101111110001010;
assign data[15][17] = 32'b00000000101000101010001010100011;
assign data[15][18] = 32'b00000000110001101100011011000111;
assign data[15][19] = 32'b00000000011010100001010011000000;
assign data[15][20] = 32'b00000000000101000110100110111111;
assign data[15][21] = 32'b00000000000000000000000000000000;
assign data[15][22] = 32'b00000000000000000000000000000000;
assign data[15][23] = 32'b00000000000000000000000000000000;
assign data[15][24] = 32'b00000000000000000000000000000000;
assign data[15][25] = 32'b00000000000000000000000000000000;
assign data[15][26] = 32'b00000000000000000000000000000000;
assign data[15][27] = 32'b00000000000000000000000000000000;
assign data[16][0] = 32'b00000000000000000000000000000000;
assign data[16][1] = 32'b00000000000000000000000000000000;
assign data[16][2] = 32'b00000000000000000000000000000000;
assign data[16][3] = 32'b00000000000000000000000000000000;
assign data[16][4] = 32'b00000000000000000000000000000000;
assign data[16][5] = 32'b00000000000000000000000000000000;
assign data[16][6] = 32'b00000000000000000000000000000000;
assign data[16][7] = 32'b00000000000000000000000000000000;
assign data[16][8] = 32'b00000000000000000000000000000000;
assign data[16][9] = 32'b00000000000000000000000000000000;
assign data[16][10] = 32'b00000000000000000000000000000000;
assign data[16][11] = 32'b00000000000000000000000000000000;
assign data[16][12] = 32'b00000000000000000000000000000000;
assign data[16][13] = 32'b00000000000000000000000000000000;
assign data[16][14] = 32'b00000000000000000000000000000000;
assign data[16][15] = 32'b00000000000100001011101101100110;
assign data[16][16] = 32'b00000000011101001100101000100000;
assign data[16][17] = 32'b00000000110011101100111011001111;
assign data[16][18] = 32'b00000000101001101010011010100111;
assign data[16][19] = 32'b00000000001101001000100111011111;
assign data[16][20] = 32'b00000000000000111010111001011001;
assign data[16][21] = 32'b00000000000000000000000000000000;
assign data[16][22] = 32'b00000000000000000000000000000000;
assign data[16][23] = 32'b00000000000000000000000000000000;
assign data[16][24] = 32'b00000000000000000000000000000000;
assign data[16][25] = 32'b00000000000000000000000000000000;
assign data[16][26] = 32'b00000000000000000000000000000000;
assign data[16][27] = 32'b00000000000000000000000000000000;
assign data[17][0] = 32'b00000000000000000000000000000000;
assign data[17][1] = 32'b00000000000000000000000000000000;
assign data[17][2] = 32'b00000000000000000000000000000000;
assign data[17][3] = 32'b00000000000000000000000000000000;
assign data[17][4] = 32'b00000000000000000000000000000000;
assign data[17][5] = 32'b00000000000000000000000000000000;
assign data[17][6] = 32'b00000000000000000000000000000000;
assign data[17][7] = 32'b00000000000000000000000000000000;
assign data[17][8] = 32'b00000000000000000000000000000000;
assign data[17][9] = 32'b00000000000000000000000000000000;
assign data[17][10] = 32'b00000000000000000000000000000000;
assign data[17][11] = 32'b00000000000000000000000000000000;
assign data[17][12] = 32'b00000000000000000000000000000000;
assign data[17][13] = 32'b00000000000000000000000000000000;
assign data[17][14] = 32'b00000000000000100000001000000010;
assign data[17][15] = 32'b00000000001110110011101100111011;
assign data[17][16] = 32'b00000000101001101111110001010010;
assign data[17][17] = 32'b00000000110000001100000011000001;
assign data[17][18] = 32'b00000000010111110101111101100000;
assign data[17][19] = 32'b00000000000100010110011010111100;
assign data[17][20] = 32'b00000000000000000101010110101011;
assign data[17][21] = 32'b00000000000000000000000000000000;
assign data[17][22] = 32'b00000000000000000000000000000000;
assign data[17][23] = 32'b00000000000000000000000000000000;
assign data[17][24] = 32'b00000000000000000000000000000000;
assign data[17][25] = 32'b00000000000000000000000000000000;
assign data[17][26] = 32'b00000000000000000000000000000000;
assign data[17][27] = 32'b00000000000000000000000000000000;
assign data[18][0] = 32'b00000000000000000000000000000000;
assign data[18][1] = 32'b00000000000000000000000000000000;
assign data[18][2] = 32'b00000000000000000000000000000000;
assign data[18][3] = 32'b00000000000000000000000000000000;
assign data[18][4] = 32'b00000000000000000000000000000000;
assign data[18][5] = 32'b00000000000000000000000000000000;
assign data[18][6] = 32'b00000000000000000000000000000000;
assign data[18][7] = 32'b00000000000000000000000000000000;
assign data[18][8] = 32'b00000000000000000000000000000000;
assign data[18][9] = 32'b00000000000000000000000000000000;
assign data[18][10] = 32'b00000000000000000000000000000000;
assign data[18][11] = 32'b00000000000000000000000000000000;
assign data[18][12] = 32'b00000000000000000000000000000000;
assign data[18][13] = 32'b00000000000000000000000000000000;
assign data[18][14] = 32'b00000000000101000001010000010100;
assign data[18][15] = 32'b00000000011101111100110100100011;
assign data[18][16] = 32'b00000000110010001100100011001001;
assign data[18][17] = 32'b00000000100101110100000111101101;
assign data[18][18] = 32'b00000000001011011101100010000011;
assign data[18][19] = 32'b00000000000000110101100010101110;
assign data[18][20] = 32'b00000000000000000000000000000000;
assign data[18][21] = 32'b00000000000000000000000000000000;
assign data[18][22] = 32'b00000000000000000000000000000000;
assign data[18][23] = 32'b00000000000000000000000000000000;
assign data[18][24] = 32'b00000000000000000000000000000000;
assign data[18][25] = 32'b00000000000000000000000000000000;
assign data[18][26] = 32'b00000000000000000000000000000000;
assign data[18][27] = 32'b00000000000000000000000000000000;
assign data[19][0] = 32'b00000000000000000000000000000000;
assign data[19][1] = 32'b00000000000000000000000000000000;
assign data[19][2] = 32'b00000000000000000000000000000000;
assign data[19][3] = 32'b00000000000000000000000000000000;
assign data[19][4] = 32'b00000000000000000000000000000000;
assign data[19][5] = 32'b00000000000000000000000000000000;
assign data[19][6] = 32'b00000000000000000000000000000000;
assign data[19][7] = 32'b00000000000000000000000000000000;
assign data[19][8] = 32'b00000000000000000000000000000000;
assign data[19][9] = 32'b00000000000000000000000000000000;
assign data[19][10] = 32'b00000000000000000000000000000000;
assign data[19][11] = 32'b00000000000000000000000000000000;
assign data[19][12] = 32'b00000000000000000000000000000000;
assign data[19][13] = 32'b00000000000000100000001000000010;
assign data[19][14] = 32'b00000000010000011110110010011000;
assign data[19][15] = 32'b00000000101100110000100001011110;
assign data[19][16] = 32'b00000000110010110010000001110110;
assign data[19][17] = 32'b00000000011001111011110100010011;
assign data[19][18] = 32'b00000000000101000001010000010100;
assign data[19][19] = 32'b00000000000000000101010110101011;
assign data[19][20] = 32'b00000000000000000000000000000000;
assign data[19][21] = 32'b00000000000000000000000000000000;
assign data[19][22] = 32'b00000000000000000000000000000000;
assign data[19][23] = 32'b00000000000000000000000000000000;
assign data[19][24] = 32'b00000000000000000000000000000000;
assign data[19][25] = 32'b00000000000000000000000000000000;
assign data[19][26] = 32'b00000000000000000000000000000000;
assign data[19][27] = 32'b00000000000000000000000000000000;
assign data[20][0] = 32'b00000000000000000000000000000000;
assign data[20][1] = 32'b00000000000000000000000000000000;
assign data[20][2] = 32'b00000000000000000000000000000000;
assign data[20][3] = 32'b00000000000000000000000000000000;
assign data[20][4] = 32'b00000000000000000000000000000000;
assign data[20][5] = 32'b00000000000000000000000000000000;
assign data[20][6] = 32'b00000000000000000000000000000000;
assign data[20][7] = 32'b00000000000000000000000000000000;
assign data[20][8] = 32'b00000000000000000000000000000000;
assign data[20][9] = 32'b00000000000000000000000000000000;
assign data[20][10] = 32'b00000000000000000000000000000000;
assign data[20][11] = 32'b00000000000000000000000000000000;
assign data[20][12] = 32'b00000000000000000000000000000000;
assign data[20][13] = 32'b00000000000100101011110101101000;
assign data[20][14] = 32'b00000000011101010001111111001011;
assign data[20][15] = 32'b00000000110011111100111111010000;
assign data[20][16] = 32'b00000000101001001010010010100101;
assign data[20][17] = 32'b00000000001100011101110010000111;
assign data[20][18] = 32'b00000000000000110000001100000011;
assign data[20][19] = 32'b00000000000000000000000000000000;
assign data[20][20] = 32'b00000000000000000000000000000000;
assign data[20][21] = 32'b00000000000000000000000000000000;
assign data[20][22] = 32'b00000000000000000000000000000000;
assign data[20][23] = 32'b00000000000000000000000000000000;
assign data[20][24] = 32'b00000000000000000000000000000000;
assign data[20][25] = 32'b00000000000000000000000000000000;
assign data[20][26] = 32'b00000000000000000000000000000000;
assign data[20][27] = 32'b00000000000000000000000000000000;
assign data[21][0] = 32'b00000000000000000000000000000000;
assign data[21][1] = 32'b00000000000000000000000000000000;
assign data[21][2] = 32'b00000000000000000000000000000000;
assign data[21][3] = 32'b00000000000000000000000000000000;
assign data[21][4] = 32'b00000000000000000000000000000000;
assign data[21][5] = 32'b00000000000000000000000000000000;
assign data[21][6] = 32'b00000000000000000000000000000000;
assign data[21][7] = 32'b00000000000000000000000000000000;
assign data[21][8] = 32'b00000000000000000000000000000000;
assign data[21][9] = 32'b00000000000000000000000000000000;
assign data[21][10] = 32'b00000000000000000000000000000000;
assign data[21][11] = 32'b00000000000000000000000000000000;
assign data[21][12] = 32'b00000000000000000000000000000000;
assign data[21][13] = 32'b00000000000110101100010101110000;
assign data[21][14] = 32'b00000000011101011100101100100001;
assign data[21][15] = 32'b00000000101101001011010010110101;
assign data[21][16] = 32'b00000000011010100110101001101011;
assign data[21][17] = 32'b00000000000101010001010100010101;
assign data[21][18] = 32'b00000000000000000000000000000000;
assign data[21][19] = 32'b00000000000000000000000000000000;
assign data[21][20] = 32'b00000000000000000000000000000000;
assign data[21][21] = 32'b00000000000000000000000000000000;
assign data[21][22] = 32'b00000000000000000000000000000000;
assign data[21][23] = 32'b00000000000000000000000000000000;
assign data[21][24] = 32'b00000000000000000000000000000000;
assign data[21][25] = 32'b00000000000000000000000000000000;
assign data[21][26] = 32'b00000000000000000000000000000000;
assign data[21][27] = 32'b00000000000000000000000000000000;
assign data[22][0] = 32'b00000000000000000000000000000000;
assign data[22][1] = 32'b00000000000000000000000000000000;
assign data[22][2] = 32'b00000000000000000000000000000000;
assign data[22][3] = 32'b00000000000000000000000000000000;
assign data[22][4] = 32'b00000000000000000000000000000000;
assign data[22][5] = 32'b00000000000000000000000000000000;
assign data[22][6] = 32'b00000000000000000000000000000000;
assign data[22][7] = 32'b00000000000000000000000000000000;
assign data[22][8] = 32'b00000000000000000000000000000000;
assign data[22][9] = 32'b00000000000000000000000000000000;
assign data[22][10] = 32'b00000000000000000000000000000000;
assign data[22][11] = 32'b00000000000000000000000000000000;
assign data[22][12] = 32'b00000000000000000000000000000000;
assign data[22][13] = 32'b00000000000010010101111010110100;
assign data[22][14] = 32'b00000000001110000011100000111000;
assign data[22][15] = 32'b00000000010101101010110000000010;
assign data[22][16] = 32'b00000000001010110010101100101011;
assign data[22][17] = 32'b00000000000001100101101110110001;
assign data[22][18] = 32'b00000000000000000000000000000000;
assign data[22][19] = 32'b00000000000000000000000000000000;
assign data[22][20] = 32'b00000000000000000000000000000000;
assign data[22][21] = 32'b00000000000000000000000000000000;
assign data[22][22] = 32'b00000000000000000000000000000000;
assign data[22][23] = 32'b00000000000000000000000000000000;
assign data[22][24] = 32'b00000000000000000000000000000000;
assign data[22][25] = 32'b00000000000000000000000000000000;
assign data[22][26] = 32'b00000000000000000000000000000000;
assign data[22][27] = 32'b00000000000000000000000000000000;
assign data[23][0] = 32'b00000000000000000000000000000000;
assign data[23][1] = 32'b00000000000000000000000000000000;
assign data[23][2] = 32'b00000000000000000000000000000000;
assign data[23][3] = 32'b00000000000000000000000000000000;
assign data[23][4] = 32'b00000000000000000000000000000000;
assign data[23][5] = 32'b00000000000000000000000000000000;
assign data[23][6] = 32'b00000000000000000000000000000000;
assign data[23][7] = 32'b00000000000000000000000000000000;
assign data[23][8] = 32'b00000000000000000000000000000000;
assign data[23][9] = 32'b00000000000000000000000000000000;
assign data[23][10] = 32'b00000000000000000000000000000000;
assign data[23][11] = 32'b00000000000000000000000000000000;
assign data[23][12] = 32'b00000000000000000000000000000000;
assign data[23][13] = 32'b00000000000000001010101101010110;
assign data[23][14] = 32'b00000000000001111011001001011101;
assign data[23][15] = 32'b00000000000011010000110100001101;
assign data[23][16] = 32'b00000000000001100000011000000110;
assign data[23][17] = 32'b00000000000000001010101101010110;
assign data[23][18] = 32'b00000000000000000000000000000000;
assign data[23][19] = 32'b00000000000000000000000000000000;
assign data[23][20] = 32'b00000000000000000000000000000000;
assign data[23][21] = 32'b00000000000000000000000000000000;
assign data[23][22] = 32'b00000000000000000000000000000000;
assign data[23][23] = 32'b00000000000000000000000000000000;
assign data[23][24] = 32'b00000000000000000000000000000000;
assign data[23][25] = 32'b00000000000000000000000000000000;
assign data[23][26] = 32'b00000000000000000000000000000000;
assign data[23][27] = 32'b00000000000000000000000000000000;
assign data[24][0] = 32'b00000000000000000000000000000000;
assign data[24][1] = 32'b00000000000000000000000000000000;
assign data[24][2] = 32'b00000000000000000000000000000000;
assign data[24][3] = 32'b00000000000000000000000000000000;
assign data[24][4] = 32'b00000000000000000000000000000000;
assign data[24][5] = 32'b00000000000000000000000000000000;
assign data[24][6] = 32'b00000000000000000000000000000000;
assign data[24][7] = 32'b00000000000000000000000000000000;
assign data[24][8] = 32'b00000000000000000000000000000000;
assign data[24][9] = 32'b00000000000000000000000000000000;
assign data[24][10] = 32'b00000000000000000000000000000000;
assign data[24][11] = 32'b00000000000000000000000000000000;
assign data[24][12] = 32'b00000000000000000000000000000000;
assign data[24][13] = 32'b00000000000000000000000000000000;
assign data[24][14] = 32'b00000000000000000000000000000000;
assign data[24][15] = 32'b00000000000000000000000000000000;
assign data[24][16] = 32'b00000000000000000000000000000000;
assign data[24][17] = 32'b00000000000000000000000000000000;
assign data[24][18] = 32'b00000000000000000000000000000000;
assign data[24][19] = 32'b00000000000000000000000000000000;
assign data[24][20] = 32'b00000000000000000000000000000000;
assign data[24][21] = 32'b00000000000000000000000000000000;
assign data[24][22] = 32'b00000000000000000000000000000000;
assign data[24][23] = 32'b00000000000000000000000000000000;
assign data[24][24] = 32'b00000000000000000000000000000000;
assign data[24][25] = 32'b00000000000000000000000000000000;
assign data[24][26] = 32'b00000000000000000000000000000000;
assign data[24][27] = 32'b00000000000000000000000000000000;
assign data[25][0] = 32'b00000000000000000000000000000000;
assign data[25][1] = 32'b00000000000000000000000000000000;
assign data[25][2] = 32'b00000000000000000000000000000000;
assign data[25][3] = 32'b00000000000000000000000000000000;
assign data[25][4] = 32'b00000000000000000000000000000000;
assign data[25][5] = 32'b00000000000000000000000000000000;
assign data[25][6] = 32'b00000000000000000000000000000000;
assign data[25][7] = 32'b00000000000000000000000000000000;
assign data[25][8] = 32'b00000000000000000000000000000000;
assign data[25][9] = 32'b00000000000000000000000000000000;
assign data[25][10] = 32'b00000000000000000000000000000000;
assign data[25][11] = 32'b00000000000000000000000000000000;
assign data[25][12] = 32'b00000000000000000000000000000000;
assign data[25][13] = 32'b00000000000000000000000000000000;
assign data[25][14] = 32'b00000000000000000000000000000000;
assign data[25][15] = 32'b00000000000000000000000000000000;
assign data[25][16] = 32'b00000000000000000000000000000000;
assign data[25][17] = 32'b00000000000000000000000000000000;
assign data[25][18] = 32'b00000000000000000000000000000000;
assign data[25][19] = 32'b00000000000000000000000000000000;
assign data[25][20] = 32'b00000000000000000000000000000000;
assign data[25][21] = 32'b00000000000000000000000000000000;
assign data[25][22] = 32'b00000000000000000000000000000000;
assign data[25][23] = 32'b00000000000000000000000000000000;
assign data[25][24] = 32'b00000000000000000000000000000000;
assign data[25][25] = 32'b00000000000000000000000000000000;
assign data[25][26] = 32'b00000000000000000000000000000000;
assign data[25][27] = 32'b00000000000000000000000000000000;
assign data[26][0] = 32'b00000000000000000000000000000000;
assign data[26][1] = 32'b00000000000000000000000000000000;
assign data[26][2] = 32'b00000000000000000000000000000000;
assign data[26][3] = 32'b00000000000000000000000000000000;
assign data[26][4] = 32'b00000000000000000000000000000000;
assign data[26][5] = 32'b00000000000000000000000000000000;
assign data[26][6] = 32'b00000000000000000000000000000000;
assign data[26][7] = 32'b00000000000000000000000000000000;
assign data[26][8] = 32'b00000000000000000000000000000000;
assign data[26][9] = 32'b00000000000000000000000000000000;
assign data[26][10] = 32'b00000000000000000000000000000000;
assign data[26][11] = 32'b00000000000000000000000000000000;
assign data[26][12] = 32'b00000000000000000000000000000000;
assign data[26][13] = 32'b00000000000000000000000000000000;
assign data[26][14] = 32'b00000000000000000000000000000000;
assign data[26][15] = 32'b00000000000000000000000000000000;
assign data[26][16] = 32'b00000000000000000000000000000000;
assign data[26][17] = 32'b00000000000000000000000000000000;
assign data[26][18] = 32'b00000000000000000000000000000000;
assign data[26][19] = 32'b00000000000000000000000000000000;
assign data[26][20] = 32'b00000000000000000000000000000000;
assign data[26][21] = 32'b00000000000000000000000000000000;
assign data[26][22] = 32'b00000000000000000000000000000000;
assign data[26][23] = 32'b00000000000000000000000000000000;
assign data[26][24] = 32'b00000000000000000000000000000000;
assign data[26][25] = 32'b00000000000000000000000000000000;
assign data[26][26] = 32'b00000000000000000000000000000000;
assign data[26][27] = 32'b00000000000000000000000000000000;
assign data[27][0] = 32'b00000000000000000000000000000000;
assign data[27][1] = 32'b00000000000000000000000000000000;
assign data[27][2] = 32'b00000000000000000000000000000000;
assign data[27][3] = 32'b00000000000000000000000000000000;
assign data[27][4] = 32'b00000000000000000000000000000000;
assign data[27][5] = 32'b00000000000000000000000000000000;
assign data[27][6] = 32'b00000000000000000000000000000000;
assign data[27][7] = 32'b00000000000000000000000000000000;
assign data[27][8] = 32'b00000000000000000000000000000000;
assign data[27][9] = 32'b00000000000000000000000000000000;
assign data[27][10] = 32'b00000000000000000000000000000000;
assign data[27][11] = 32'b00000000000000000000000000000000;
assign data[27][12] = 32'b00000000000000000000000000000000;
assign data[27][13] = 32'b00000000000000000000000000000000;
assign data[27][14] = 32'b00000000000000000000000000000000;
assign data[27][15] = 32'b00000000000000000000000000000000;
assign data[27][16] = 32'b00000000000000000000000000000000;
assign data[27][17] = 32'b00000000000000000000000000000000;
assign data[27][18] = 32'b00000000000000000000000000000000;
assign data[27][19] = 32'b00000000000000000000000000000000;
assign data[27][20] = 32'b00000000000000000000000000000000;
assign data[27][21] = 32'b00000000000000000000000000000000;
assign data[27][22] = 32'b00000000000000000000000000000000;
assign data[27][23] = 32'b00000000000000000000000000000000;
assign data[27][24] = 32'b00000000000000000000000000000000;
assign data[27][25] = 32'b00000000000000000000000000000000;
assign data[27][26] = 32'b00000000000000000000000000000000;
assign data[27][27] = 32'b00000000000000000000000000000000;


	always @(*) begin
		if (data_read_done == 1'b0) begin
			// row 0
			data_00 = data[count_x][count_y];
			data_01 = data[count_x][count_y+1];
			data_02 = data[count_x][count_y+2];
			data_03 = data[count_x][count_y+3];
			data_04 = data[count_x][count_y+4];
			// row 1
			data_10 = data[count_x+1][count_y];
			data_11 = data[count_x+1][count_y+1];
			data_12 = data[count_x+1][count_y+2];
			data_13 = data[count_x+1][count_y+3];
			data_14 = data[count_x+1][count_y+4];
			// row 2
			data_20 = data[count_x+2][count_y];
			data_21 = data[count_x+2][count_y+1];
			data_22 = data[count_x+2][count_y+2];
			data_23 = data[count_x+2][count_y+3];
			data_24 = data[count_x+2][count_y+4];
			// row 3
			data_30 = data[count_x+3][count_y];
			data_31 = data[count_x+3][count_y+1];
			data_32 = data[count_x+3][count_y+2];
			data_33 = data[count_x+3][count_y+3];
			data_34 = data[count_x+3][count_y+4];
			// row 4
			data_40 = data[count_x+4][count_y];
			data_41 = data[count_x+4][count_y+1];
			data_42 = data[count_x+4][count_y+2];
			data_43 = data[count_x+4][count_y+3];
			data_44 = data[count_x+4][count_y+4];
		end
	end

	always @(*) begin
		// depth 0
		pool_0_00 = relu_1[2*relu_count_x][2*relu_count_y];
		pool_0_01 = relu_1[2*relu_count_x][2*relu_count_y+1];
		pool_0_10 = relu_1[2*relu_count_x+1][2*relu_count_y];
		pool_0_11 = relu_1[2*relu_count_x+1][2*relu_count_y+1];
		// depth 1
		pool_1_00 = relu_2[2*relu_count_x][2*relu_count_y];
		pool_1_01 = relu_2[2*relu_count_x][2*relu_count_y+1];
		pool_1_10 = relu_2[2*relu_count_x+1][2*relu_count_y];
		pool_1_11 = relu_2[2*relu_count_x+1][2*relu_count_y+1];
		// depth 2
		pool_2_00 = relu_3[2*relu_count_x][2*relu_count_y];
		pool_2_01 = relu_3[2*relu_count_x][2*relu_count_y+1];
		pool_2_10 = relu_3[2*relu_count_x+1][2*relu_count_y];
		pool_2_11 = relu_3[2*relu_count_x+1][2*relu_count_y+1];
		// depth 3
		pool_3_00 = relu_4[2*relu_count_x][2*relu_count_y];
		pool_3_01 = relu_4[2*relu_count_x][2*relu_count_y+1];
		pool_3_10 = relu_4[2*relu_count_x+1][2*relu_count_y];
		pool_3_11 = relu_4[2*relu_count_x+1][2*relu_count_y+1];
		// depth 4
		pool_4_00 = relu_5[2*relu_count_x][2*relu_count_y];
		pool_4_01 = relu_5[2*relu_count_x][2*relu_count_y+1];
		pool_4_10 = relu_5[2*relu_count_x+1][2*relu_count_y];
		pool_4_11 = relu_5[2*relu_count_x+1][2*relu_count_y+1];
		// depth 5
		pool_5_00 = relu_6[2*relu_count_x][2*relu_count_y];
		pool_5_01 = relu_6[2*relu_count_x][2*relu_count_y+1];
		pool_5_10 = relu_6[2*relu_count_x+1][2*relu_count_y];
		pool_5_11 = relu_6[2*relu_count_x+1][2*relu_count_y+1];
		// depth 6
		pool_6_00 = relu_7[2*relu_count_x][2*relu_count_y];
		pool_6_01 = relu_7[2*relu_count_x][2*relu_count_y+1];
		pool_6_10 = relu_7[2*relu_count_x+1][2*relu_count_y];
		pool_6_11 = relu_7[2*relu_count_x+1][2*relu_count_y+1];
		// depth 7
		pool_7_00 = relu_8[2*relu_count_x][2*relu_count_y];
		pool_7_01 = relu_8[2*relu_count_x][2*relu_count_y+1];
		pool_7_10 = relu_8[2*relu_count_x+1][2*relu_count_y];
		pool_7_11 = relu_8[2*relu_count_x+1][2*relu_count_y+1];
	end

	always @(posedge clk) begin
		if (rst) count <= 0;
		else count = count + 1;
	end

	always @(posedge clk) begin
		if (rst) begin
			count_x <= 0;
			count_y <= 0;
		end else if (count_y < 5'd23) begin
			count_y <= count_y + 1;
		end else if (count_y == 5'd23) begin
			count_x <= count_x + 1;
			count_y <= 0;
		end

		if (rst) begin
			data_read_done <= 1'b0;
		end else if (count_y == 5'd23 && count_x == 5'd23) begin
			data_read_done <= 1'b1;
		end
	end

	always @(posedge clk) begin
		if (rst) begin
			relu_count_x <= 0;
			relu_count_y <= 0;
		end else if (count >=579 && count < 723) begin
			if (relu_count_y < 5'd11) begin
				relu_count_y <= relu_count_y + 1;
			end else if (relu_count_y == 5'd11) begin
				relu_count_x <= relu_count_x + 1;
				relu_count_y <= 0;
			end
		end
	end

	always @(*) begin
		if (count > 1 && count <578) begin
			relu[0][count-2] = relu_result_1;
			relu[1][count-2] = relu_result_2;
			relu[2][count-2] = relu_result_3;
			relu[3][count-2] = relu_result_4;
			relu[4][count-2] = relu_result_5;
			relu[5][count-2] = relu_result_6;
			relu[6][count-2] = relu_result_7;
			relu[7][count-2] = relu_result_8;
		end
	end

	always @(*) begin
		for (i = 0; i < 24; i = i+1) begin
			for (j = 0; j < 24; j = j+1) begin
				relu_1[i][j] = relu[0][24*i + j];
				relu_2[i][j] = relu[1][24*i + j];
				relu_3[i][j] = relu[2][24*i + j];
				relu_4[i][j] = relu[3][24*i + j];
				relu_5[i][j] = relu[4][24*i + j];
				relu_6[i][j] = relu[5][24*i + j];
				relu_7[i][j] = relu[6][24*i + j];
				relu_8[i][j] = relu[7][24*i + j];
			end
		end
	end

	conv_layer conv(
		// INPUTS
	 	.clk(clk),
	 	.rst(rst),
		.data_00(data_00),
		.data_01(data_01),
		.data_02(data_02),
		.data_03(data_03),
		.data_04(data_04),
		.data_10(data_10),
		.data_11(data_11),
		.data_12(data_12),
		.data_13(data_13),
		.data_14(data_14),
		.data_20(data_20),
		.data_21(data_21),
		.data_22(data_22),
		.data_23(data_23),
		.data_24(data_24),
		.data_30(data_30),
		.data_31(data_31),
		.data_32(data_32),
		.data_33(data_33),
		.data_34(data_34),
		.data_40(data_40),
		.data_41(data_41),
		.data_42(data_42),
		.data_43(data_43),
		.data_44(data_44),
		// OUTPUTS
	 	.conv_result_1(conv_result_1),
	 	.conv_result_2(conv_result_2),
	 	.conv_result_3(conv_result_3),
	 	.conv_result_4(conv_result_4),
	 	.conv_result_5(conv_result_5),
	 	.conv_result_6(conv_result_6),
	 	.conv_result_7(conv_result_7),
	 	.conv_result_8(conv_result_8)
	);

	relu_layer relu_l(
		// INPUTS
		.clk(clk),
	 	.rst(rst),
		.conv_result_1(conv_result_1),
		.conv_result_2(conv_result_2),
		.conv_result_3(conv_result_3),
		.conv_result_4(conv_result_4),
		.conv_result_5(conv_result_5),
		.conv_result_6(conv_result_6),
		.conv_result_7(conv_result_7),
		.conv_result_8(conv_result_8),
		// OUTPUTS
		.relu_result_1(relu_result_1),
		.relu_result_2(relu_result_2),
		.relu_result_3(relu_result_3),
		.relu_result_4(relu_result_4),
		.relu_result_5(relu_result_5),
		.relu_result_6(relu_result_6),
		.relu_result_7(relu_result_7),
		.relu_result_8(relu_result_8)
	);

// pool_layer
	pool_layer pool_l(
		// INPUTS
		.clk(clk),
	 	.rst(rst),
		.count_x(relu_count_x),
		.count_y(relu_count_y),
		.pool_0_00 (pool_0_00),
		.pool_0_01 (pool_0_01),
		.pool_0_10 (pool_0_10),
		.pool_0_11 (pool_0_11),
		.pool_1_00 (pool_1_00),
		.pool_1_01 (pool_1_01),
		.pool_1_10 (pool_1_10),
		.pool_1_11 (pool_1_11),
		.pool_2_00 (pool_2_00),
		.pool_2_01 (pool_2_01),
		.pool_2_10 (pool_2_10),
		.pool_2_11 (pool_2_11),
		.pool_3_00 (pool_3_00),
		.pool_3_01 (pool_3_01),
		.pool_3_10 (pool_3_10),
		.pool_3_11 (pool_3_11),
		.pool_4_00 (pool_4_00),
		.pool_4_01 (pool_4_01),
		.pool_4_10 (pool_4_10),
		.pool_4_11 (pool_4_11),
		.pool_5_00 (pool_5_00),
		.pool_5_01 (pool_5_01),
		.pool_5_10 (pool_5_10),
		.pool_5_11 (pool_5_11),
		.pool_6_00 (pool_6_00),
		.pool_6_01 (pool_6_01),
		.pool_6_10 (pool_6_10),
		.pool_6_11 (pool_6_11),
		.pool_7_00 (pool_7_00),
		.pool_7_01 (pool_7_01),
		.pool_7_10 (pool_7_10),
		.pool_7_11 (pool_7_11),
		// OUTPUTS
		/*
		.pool_result_1(pool_result_1),
		.pool_result_2(pool_result_2),
		.pool_result_3(pool_result_3),
		.pool_result_4(pool_result_4),
		.pool_result_5(pool_result_5),
		.pool_result_6(pool_result_6),
		.pool_result_7(pool_result_7),
		.pool_result_8(pool_result_8)
		*/
		.prob_0(prob_0),
		.prob_1(prob_1),
		.prob_2(prob_2),
		.prob_3(prob_3),
		.prob_4(prob_4),
		.prob_5(prob_5),
		.prob_6(prob_6),
		.prob_7(prob_7),
		.prob_8(prob_8),
		.prob_9(prob_9),
		.fc_done(fc_done)
	);
	/*
	// fc_layer
		fc_layer fc(
			// INPUTS
			.clk(clk),
		 	.rst(rst),
			.fc_enable(pool_done),
			.pool_result_1(pool_result_1),
			.pool_result_2(pool_result_2),
			.pool_result_3(pool_result_3),
			.pool_result_4(pool_result_4),
			.pool_result_5(pool_result_5),
			.pool_result_6(pool_result_6),
			.pool_result_7(pool_result_7),
			.pool_result_8(pool_result_8),
			.fc_weight_0(fc_weight_0),
			.fc_weight_1(fc_weight_1),
			.fc_weight_2(fc_weight_2),
			.fc_weight_3(fc_weight_3),
			.fc_weight_4(fc_weight_4),
			.fc_weight_5(fc_weight_5),
			.fc_weight_6(fc_weight_6),
			.fc_weight_7(fc_weight_7),
			.fc_weight_8(fc_weight_8),
			.fc_weight_9(fc_weight_9),

			// OUTPUTS
			.prob_0(prob_0),
			.prob_1(prob_1),
			.prob_2(prob_2),
			.prob_3(prob_3),
			.prob_4(prob_4),
			.prob_5(prob_5),
			.prob_6(prob_6),
			.prob_7(prob_7),
			.prob_8(prob_8),
			.prob_9(prob_9),
			.fc_done(fc_done)
		);
		*/
// Compare prob0-prob9 and get result

	reg signed [112:0] in_prob_0, in_prob_1, in_prob_2, in_prob_3, in_prob_4, in_prob_5, in_prob_6, in_prob_7, in_prob_8, in_prob_9;

	always @ (fc_done) begin
		in_prob_0 = prob_0;
		in_prob_1 = prob_1;
		in_prob_2 = prob_2;
		in_prob_3 = prob_3;
		in_prob_4 = prob_4;
		in_prob_5 = prob_5;
		in_prob_6 = prob_6;
		in_prob_7 = prob_7;
		in_prob_8 = prob_8;
		in_prob_9 = prob_9;
	end

	reg signed [112:0] tmp_prob;
	reg [3:0] next_result;
	reg signed [112:0] max_prob;

	always @ (*) begin
		prob[0] = in_prob_0;
		prob[1] = in_prob_1;
		prob[2] = in_prob_2;
		prob[3] = in_prob_3;
		prob[4] = in_prob_4;
		prob[5] = in_prob_5;
		prob[6] = in_prob_6;
		prob[7] = in_prob_7;
		prob[8] = in_prob_8;
		prob[9] = in_prob_9;
		next_result = 0;
		max_prob = prob[0];
		for (i = 1; i < 10; i=i+1) begin
			if (max_prob < prob[i]) begin
				max_prob = prob[i];
				next_result = i;
			end
		end
	end

	always @ (posedge clk) begin
		if (rst) result <= 0;
		else result <= next_result;
	end
endmodule
